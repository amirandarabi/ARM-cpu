module CPU();
clock c(clk);
endmodule 