module RUN();
clock c(clk);
testbench tb(clk);
endmodule 